$date
   Sun Mar 23 19:26:55 2025
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module serial_tb $end
$var wire 1 ! uart_line $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
1!
$end
#13150000
0!
#48990000
1!
#57950000
0!
#66910000
1!
#75870000
0!
#84830000
1!
#93790000
0!
#102750000
1!
#147550000
0!
#156510000
1!
#165470000
0!
#174430000
1!
#210270000
0!
#219230000
1!
#281950000
0!
#290910000
1!
#317790000
0!
#326750000
1!
#335710000
0!
#362590000
1!
#416350000
0!
#470110000
1!
#496990000
0!
#505950000
1!
#550750000
0!
#568670000
1!
#577630000
0!
#613470000
1!
#631390000
0!
#640350000
1!
#685150000
0!
#694110000
1!
#712030000
0!
#765790000
1!
#819550000
0!
#828510000
1!
#953950000
0!
#971870000
1!
#989790000
0!
#1016670000
1!
#1025630000
0!
#1043550000
1!
