$date
   Sat Mar  8 13:06:12 2025
$end
$version
  2023.1
$end
$timescale
  1ps
$end
$scope module Sequence_Detector_tb $end
$var wire 1 " reset $end
$var wire 1 ! clock $end
$var wire 1 # load $end
$var wire 16 & input $end
$var wire 1 $ Y $end
$var wire 1 % shift_left $end
$var wire 16 ' output_structural $end
$var wire 16 -! output_behavioral $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
bx !!
1"
b0 "!
0#
x#!
0$
bx0 $!
0%
x%!
b0 &
x&!
bx '
bx '!
bx (
b0 (!
bx )
x)!
bx *
bx0 *!
bx +
x+!
b0 ,
x,!
x-
b0 -!
bx0 .
b0 .!
x/
x0
bx 1
b0 2
x3
bx0 4
x5
x6
bx 7
b0 8
x9
bx0 :
x;
x<
bx =
b0 >
x?
bx0 @
xA
xB
bx C
b0 D
xE
bx0 F
xG
xH
bx I
b0 J
xK
bx0 L
xM
xN
bx O
b0 P
xQ
bx0 R
xS
xT
bx U
b0 V
xW
bx0 X
xY
xZ
bx [
b0 \
x]
bx0 ^
x_
x`
bx a
b0 b
xc
bx0 d
xe
xf
bx g
b0 h
xi
bx0 j
xk
xl
bx m
b0 n
xo
bx0 p
xq
xr
bx s
b0 t
xu
bx0 v
xw
xx
bx y
b0 z
x{
bx0 |
x}
x~
$end
#5000
1!
b0 '
b0 (
b0 )
b0 *
b0 1
06
0c
0e
0f
#10000
0!
#15000
1!
#20000
0!
#25000
1!
#30000
0!
#35000
1!
#40000
0!
#45000
1!
#50000
0!
#55000
1!
#60000
0!
#65000
1!
#70000
0!
#75000
1!
#80000
0!
#85000
1!
#90000
0!
#95000
1!
#100000
0!
0"
1#
b0 $!
b110111101011101 &
b110111101011101 *
1+!
b0 .
b1 4
15
b1 :
1;
b0 @
1G
b1 L
1M
1S
b1 X
1Y
b0 ^
b1 d
1e
b0 j
b1 p
1q
1w
1}
#105000
1!
b1110 !!
1#!
b10 $!
b110111101011101 '
b101 '!
b110111101011101 (
b1011011110101110 )
b1011 +
1,!
1-
b110111101011101 -!
b10 .
b110111101011101 .!
b110 1
16
b1001 7
19
b11 :
1<
b1111 =
1?
b10 @
b111 C
1H
b1011 I
1K
b11 L
1N
b1110 O
1Q
b11 R
1T
b1101 U
1W
b11 X
1Z
b1110 [
1]
b10 ^
b101 a
1f
b1011 g
1i
b10 j
b111 m
1r
b1010 s
1u
b11 v
1x
b1101 y
1{
b11 |
1~
#110000
0!
0#
1%!
b1011011110101110 *
1/
05
1A
1_
0e
1k
#115000
1!
b1101 !!
1&!
b1011011110101110 '
b1110 '!
b1011011110101110 (
b101101111010111 )
1)!
b101101111010111 *
b11 *!
b101 +
1+!
0-
b1011011110101110 -!
b0 .
b1011011110101110 .!
0/
10
b1011 1
13
b11 4
15
06
b110 7
b1 :
b1001 =
1B
b1111 C
1E
b11 F
1G
b111 I
b1 L
b1011 O
b1110 U
b1101 [
1`
b1110 a
1c
b11 d
1e
0f
b101 g
b0 j
1l
b1011 m
1o
b11 p
1q
b111 s
b1 v
b1010 y
#120000
0!
b10 "!
b0 $!
1%
b10 (!
b110111101011101 )
b110111101011101 *
b10 ,
b10 2
b10 8
19
b11 :
1;
b10 >
b0 @
b10 D
b10 J
1K
b11 L
1M
b10 P
b10 V
b10 \
0]
b0 ^
0_
b10 b
b10 h
b10 n
b10 t
1u
b11 v
1w
b10 z
#125000
1!
b1110 !!
1#!
b10 $!
1%!
b110111101011101 '
b101 '!
b110111101011101 (
b1101111010111010 )
b1101111010111010 *
b1 *!
b1011 +
1,!
1-
b110111101011101 -!
b10 .
b110111101011101 .!
1/
00
b110 1
16
b1001 7
b1 :
b1111 =
1?
b10 @
1A
b111 C
1H
b1011 I
b1101 U
b1 X
b1110 [
1]
b10 ^
1_
0`
b101 a
0c
b1 d
0e
1f
b1011 g
1i
b10 j
1k
b111 m
1r
b1010 s
b1101 y
b1 |
#130000
0!
1$
b0 $!
b1011110101110101 )
1)!
b1011110101110101 *
b11 *!
1+!
03
b1 4
05
19
b11 :
1;
b1 R
1W
b11 X
1Y
0]
b0 ^
0_
1c
b11 d
1e
b1 v
1{
b11 |
1}
#135000
1!
b1011 !!
1#!
b10 $!
1%!
b1011110101110101 '
b110 '!
b1011110101110101 (
b1111010111010110 )
b1111010111010110 *
b1 *!
b1011110101110101 -!
b1011110101110101 .!
10
b1111 1
13
b11 4
15
06
b111 7
b1011 =
1B
b1110 C
b1 F
b101 U
b1011 [
1]
b10 ^
1_
b111 a
b0 j
1l
b1101 m
b101 y
#140000
0!
b1 "!
b0 $!
0%
b1 (!
b110111101011101 )
1)!
b110111101011101 *
b11 *!
1+!
b1 ,
0-
b0 .
0/
b1 2
b1 8
b1 >
b0 @
b1 D
1E
b11 F
1G
b1 J
b1 P
1Q
b11 R
1S
b1 V
b1 \
0]
b0 ^
0_
b1 b
b1 h
b1 n
b1 t
1u
b11 v
1w
b1 z
#145000
1!
1#!
b10 $!
1%!
b110111101011101 '
b101 '!
b110111101011101 (
b101101111010111 )
b101101111010111 *
b1011 +
b110111101011101 -!
b110111101011101 .!
00
b110 1
16
b1001 7
b1 :
1?
b10 @
1A
b111 C
b1011 I
b1 L
1T
b1101 U
b10 ^
b1011 g
b111 m
b1010 s
b1 v
1x
b1101 y
